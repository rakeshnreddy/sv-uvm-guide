`define uvm_object_utils(x)
`define uvm_component_utils(x)
