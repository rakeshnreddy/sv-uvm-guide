package uvm_pkg;
  class uvm_object; endclass
  class uvm_component; endclass
  class uvm_reg; endclass
  class uvm_reg_field; endclass
  class uvm_reg_block; endclass
  class uvm_sequence_item; endclass
  class uvm_sequence #(type T=int); endclass
  class uvm_sequencer #(type T=int); endclass
  class uvm_phase; endclass
  class uvm_reg_item; endclass
  class uvm_reg_predictor; endclass
  typedef int uvm_status_e;
endpackage
