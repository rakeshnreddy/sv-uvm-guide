`ifndef SEQUENCER_SV
`define SEQUENCER_SV

typedef uvm_sequencer #(sequence_item) sequencer;

`endif // SEQUENCER_SV
